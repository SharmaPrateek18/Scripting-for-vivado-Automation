module top_CLA16(output [15:0] sum, output cout, input [15:0] a, b);
wire [2079:0] g, p, c;
wire [135:0] e;
wire cin;
buf #(1) (cin, 0);
//c[0]
and #(1) (e[0], cin, p[0]);
or #(1) (c[0], e[0], g[0]);

//c[1]
and #(1) (e[1], cin, p[0], p[1]);
and #(1) (e[2], g[0], p[1]);
or #(1) (c[1], e[1], e[2], g[1]);

//c[2]
and #(1) (e[3], cin, p[0], p[1], p[2]);
and #(1) (e[4], g[0], p[1], p[2]);
and #(1) (e[5], g[1], p[2]);
or #(1) (c[2], e[3], e[4], e[5], g[2]);

//c[3]
and #(1) (e[6], cin, p[0], p[1], p[2], p[3]);
and #(1) (e[7], g[0], p[1], p[2], p[3]);
and #(1) (e[8], g[1], p[2], p[3]);
and #(1) (e[9], g[2], p[3]);
or #(1) (c[3], e[6], e[7], e[8], e[9], g[3]);

//c[4]
and #(1) (e[10], cin, p[0], p[1], p[2], p[3], p[4]);
and #(1) (e[11], g[0], p[1], p[2], p[3], p[4]);
and #(1) (e[12], g[1], p[2], p[3], p[4]);
and #(1) (e[13], g[2], p[3], p[4]);
and #(1) (e[14], g[3], p[4]);
or #(1) (c[4], e[10], e[11], e[12], e[13], e[14], g[4]);

//c[5]
and #(1) (e[15], cin, p[0], p[1], p[2], p[3], p[4], p[5]);
and #(1) (e[16], g[0], p[1], p[2], p[3], p[4], p[5]);
and #(1) (e[17], g[1], p[2], p[3], p[4], p[5]);
and #(1) (e[18], g[2], p[3], p[4], p[5]);
and #(1) (e[19], g[3], p[4], p[5]);
and #(1) (e[20], g[4], p[5]);
or #(1) (c[5], e[15], e[16], e[17], e[18], e[19], e[20], g[5]);

//c[6]
and #(1) (e[21], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6]);
and #(1) (e[22], g[0], p[1], p[2], p[3], p[4], p[5], p[6]);
and #(1) (e[23], g[1], p[2], p[3], p[4], p[5], p[6]);
and #(1) (e[24], g[2], p[3], p[4], p[5], p[6]);
and #(1) (e[25], g[3], p[4], p[5], p[6]);
and #(1) (e[26], g[4], p[5], p[6]);
and #(1) (e[27], g[5], p[6]);
or #(1) (c[6], e[21], e[22], e[23], e[24], e[25], e[26], e[27], g[6]);

//c[7]
and #(1) (e[28], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7]);
and #(1) (e[29], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7]);
and #(1) (e[30], g[1], p[2], p[3], p[4], p[5], p[6], p[7]);
and #(1) (e[31], g[2], p[3], p[4], p[5], p[6], p[7]);
and #(1) (e[32], g[3], p[4], p[5], p[6], p[7]);
and #(1) (e[33], g[4], p[5], p[6], p[7]);
and #(1) (e[34], g[5], p[6], p[7]);
and #(1) (e[35], g[6], p[7]);
or #(1) (c[7], e[28], e[29], e[30], e[31], e[32], e[33], e[34], e[35], g[7]);

//c[8]
and #(1) (e[36], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8]);
and #(1) (e[37], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8]);
and #(1) (e[38], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8]);
and #(1) (e[39], g[2], p[3], p[4], p[5], p[6], p[7], p[8]);
and #(1) (e[40], g[3], p[4], p[5], p[6], p[7], p[8]);
and #(1) (e[41], g[4], p[5], p[6], p[7], p[8]);
and #(1) (e[42], g[5], p[6], p[7], p[8]);
and #(1) (e[43], g[6], p[7], p[8]);
and #(1) (e[44], g[7], p[8]);
or #(1) (c[8], e[36], e[37], e[38], e[39], e[40], e[41], e[42], e[43], e[44], g[8]);

//c[9]
and #(1) (e[45], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9]);
and #(1) (e[46], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9]);
and #(1) (e[47], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9]);
and #(1) (e[48], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9]);
and #(1) (e[49], g[3], p[4], p[5], p[6], p[7], p[8], p[9]);
and #(1) (e[50], g[4], p[5], p[6], p[7], p[8], p[9]);
and #(1) (e[51], g[5], p[6], p[7], p[8], p[9]);
and #(1) (e[52], g[6], p[7], p[8], p[9]);
and #(1) (e[53], g[7], p[8], p[9]);
and #(1) (e[54], g[8], p[9]);
or #(1) (c[9], e[45], e[46], e[47], e[48], e[49], e[50], e[51], e[52], e[53], e[54], g[9]);

//c[10]
and #(1) (e[55], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10]);
and #(1) (e[56], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10]);
and #(1) (e[57], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10]);
and #(1) (e[58], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10]);
and #(1) (e[59], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10]);
and #(1) (e[60], g[4], p[5], p[6], p[7], p[8], p[9], p[10]);
and #(1) (e[61], g[5], p[6], p[7], p[8], p[9], p[10]);
and #(1) (e[62], g[6], p[7], p[8], p[9], p[10]);
and #(1) (e[63], g[7], p[8], p[9], p[10]);
and #(1) (e[64], g[8], p[9], p[10]);
and #(1) (e[65], g[9], p[10]);
or #(1) (c[10], e[55], e[56], e[57], e[58], e[59], e[60], e[61], e[62], e[63], e[64], e[65], g[10]);

//c[11]
and #(1) (e[66], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11]);
and #(1) (e[67], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11]);
and #(1) (e[68], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11]);
and #(1) (e[69], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11]);
and #(1) (e[70], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11]);
and #(1) (e[71], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11]);
and #(1) (e[72], g[5], p[6], p[7], p[8], p[9], p[10], p[11]);
and #(1) (e[73], g[6], p[7], p[8], p[9], p[10], p[11]);
and #(1) (e[74], g[7], p[8], p[9], p[10], p[11]);
and #(1) (e[75], g[8], p[9], p[10], p[11]);
and #(1) (e[76], g[9], p[10], p[11]);
and #(1) (e[77], g[10], p[11]);
or #(1) (c[11], e[66], e[67], e[68], e[69], e[70], e[71], e[72], e[73], e[74], e[75], e[76], e[77], g[11]);

//c[12]
and #(1) (e[78], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12]);
and #(1) (e[79], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12]);
and #(1) (e[80], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12]);
and #(1) (e[81], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12]);
and #(1) (e[82], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12]);
and #(1) (e[83], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12]);
and #(1) (e[84], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12]);
and #(1) (e[85], g[6], p[7], p[8], p[9], p[10], p[11], p[12]);
and #(1) (e[86], g[7], p[8], p[9], p[10], p[11], p[12]);
and #(1) (e[87], g[8], p[9], p[10], p[11], p[12]);
and #(1) (e[88], g[9], p[10], p[11], p[12]);
and #(1) (e[89], g[10], p[11], p[12]);
and #(1) (e[90], g[11], p[12]);
or #(1) (c[12], e[78], e[79], e[80], e[81], e[82], e[83], e[84], e[85], e[86], e[87], e[88], e[89], e[90], g[12]);

//c[13]
and #(1) (e[91], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[92], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[93], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[94], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[95], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[96], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[97], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[98], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[99], g[7], p[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[100], g[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[101], g[9], p[10], p[11], p[12], p[13]);
and #(1) (e[102], g[10], p[11], p[12], p[13]);
and #(1) (e[103], g[11], p[12], p[13]);
and #(1) (e[104], g[12], p[13]);
or #(1) (c[13], e[91], e[92], e[93], e[94], e[95], e[96], e[97], e[98], e[99], e[100], e[101], e[102], e[103], e[104], g[13]);

//c[14]
and #(1) (e[105], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[106], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[107], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[108], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[109], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[110], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[111], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[112], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[113], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[114], g[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[115], g[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[116], g[10], p[11], p[12], p[13], p[14]);
and #(1) (e[117], g[11], p[12], p[13], p[14]);
and #(1) (e[118], g[12], p[13], p[14]);
and #(1) (e[119], g[13], p[14]);
or #(1) (c[14], e[105], e[106], e[107], e[108], e[109], e[110], e[111], e[112], e[113], e[114], e[115], e[116], e[117], e[118], e[119], g[14]);

//c[15]
and #(1) (e[120], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[121], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[122], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[123], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[124], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[125], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[126], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[127], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[128], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[129], g[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[130], g[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[131], g[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[132], g[11], p[12], p[13], p[14], p[15]);
and #(1) (e[133], g[12], p[13], p[14], p[15]);
and #(1) (e[134], g[13], p[14], p[15]);
and #(1) (e[135], g[14], p[15]);
or #(1) (c[15], e[120], e[121], e[122], e[123], e[124], e[125], e[126], e[127], e[128], e[129], e[130], e[131], e[132], e[133], e[134], e[135], g[15]);

xor #(2) (sum[0],p[0],cin);
xor #(2) x[15:1](sum[15:1],p[15:1],c[14:0]);
buf #(1) (cout, c[15]);
PGGen pggen[15:0](g[15:0],p[15:0],a[15:0],b[15:0]);
 
endmodule
